`timescale 1ns / 1ps

module InstructionMemory (
    input [31:0] read_addr,
    output wire [31:0] instruction
);
    
    // set a size for the instruction memory
    reg[31:0] mem[49:0];
    initial begin 
        mem[0] = 32'b00100000000010000000000000100000;
        mem[1] = 32'b00100000000010010000000000110111;
        mem[2] = 32'b00000001000010011000000000100100;
        mem[3] = 32'b00000001000010011000000000100101;
        mem[4] = 32'b10101100000100000000000000000100;
        mem[5] = 32'b10101100000010000000000000001000;
        mem[6] = 32'b00000001000010011000100000100000;
        mem[7] = 32'b00000001000010011001000000100010;
        mem[8] = 32'b00100000000010000000000000100000;
        mem[9] = 32'b00100000000010000000000000100000;
        mem[10] = 32'b00100000000010000000000000100000;
        mem[11] = 32'b00010010001100100000000000010010;
        mem[12] = 32'b10001100000100010000000000000100;
        mem[13] = 32'b00110010001100100000000001001000;
        mem[14] = 32'b00100000000010000000000000100000;
        mem[15] = 32'b00100000000010000000000000100000;
        mem[16] = 32'b00100000000010000000000000100000;
        mem[17] = 32'b00010010001100100000000000001111;
        mem[18] = 32'b10001100000100110000000000001000;
        mem[19] = 32'b00100000000010000000000000100000;
        mem[20] = 32'b00100000000010000000000000100000;
        mem[21] = 32'b00100000000010000000000000100000;
        mem[22] = 32'b00010010000100110000000000001101;
        mem[23] = 32'b00000010010100011010000000101010;
        mem[24] = 32'b00100000000010000000000000100000;
        mem[25] = 32'b00100000000010000000000000100000;
        mem[26] = 32'b00100000000010000000000000100000;
        mem[27] = 32'b00010010100000000000000000001111;
        mem[28] = 32'b00000010001000001001000000100000;
        mem[29] = 32'b00001000000000000000000000010111;
        mem[30] = 32'b00100000000010000000000000000000;
        mem[31] = 32'b00100000000010010000000000000000;
        mem[32] = 32'b00001000000000000000000000111111;
        mem[33] = 32'b00100000000010000000000000000001;
        mem[34] = 32'b00100000000010010000000000000001;
        mem[35] = 32'b00001000000000000000000000111111;
        mem[36] = 32'b00100000000010000000000000000010;
        mem[37] = 32'b00100000000010010000000000000010;
        mem[38] = 32'b00001000000000000000000000111111;
        mem[39] = 32'b00100000000010000000000000000011;
        mem[40] = 32'b00100000000010010000000000000011;
        mem[41] = 32'b00001000000000000000000000111111;
    end
    
    assign instruction = mem[read_addr >> 2];

endmodule